module instructionfetch
(
);

endmodule
