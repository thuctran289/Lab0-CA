module testmux2to1
();
endmodule